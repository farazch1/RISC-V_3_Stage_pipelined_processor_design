module mux_2x1(

    );
endmodule
